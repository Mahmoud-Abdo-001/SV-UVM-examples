package shared_pkg;

parameter DATA_WIDTH = 32;
parameter ADDR_WIDTH = 8;

parameter clkprd = 10;

endpackage